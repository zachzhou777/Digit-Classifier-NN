/* Weighted binary stochastic number generator as proposed by Gupta and Kumaresan. For a schematic of 
 * the intended circuit, refer to the Survey of Stochastic Computing paper, specifically Fig. 5. */
module weighted_binary_generator(binary_number, random_number, stochastic_number);

// 'binary_number' is equivalent to the real number in the range [0,1] that the stochastic number 
// represents multiplied by 1,024. 'random_number' is a random 10-bit number such that each possible 
// 10-bit number has equal likelihood of being the value of 'random_number'
input [9:0] binary_number, random_number;

// 'stochastic_number' is the current bit being generated by the bitstream
output stochastic_number;

// 'weights' and 'intermediates' are intermediate values used in the assignment of 'stochastic_number'; 
// when referring to Fig. 5 from the Survey of Stochastic Computing paper, 'weights' correspond to Wi, 
// and 'intermediates' are the unlabeled inputs to the OR gate
wire [9:0] weights, intermediates;

// Loop counter
genvar i;

// Assign values for the weights
assign weights[9] = random_number[9];
assign weights[8] = ~random_number[9] & random_number[8];
assign weights[7] = ~random_number[9] & ~random_number[8] & random_number[7];
assign weights[6] = ~random_number[9] & ~random_number[8] & ~random_number[7] & random_number[6];
assign weights[5] = ~random_number[9] & ~random_number[8] & ~random_number[7] & ~random_number[6] & 
				random_number[5];
assign weights[4] = ~random_number[9] & ~random_number[8] & ~random_number[7] & ~random_number[6] & 
				~random_number[5] & random_number[4];
assign weights[3] = ~random_number[9] & ~random_number[8] & ~random_number[7] & ~random_number[6] & 
				~random_number[5] & ~random_number[4] & random_number[3];
assign weights[2] = ~random_number[9] & ~random_number[8] & ~random_number[7] & ~random_number[6] & 
				~random_number[5] & ~random_number[4] & ~random_number[3] & 
				random_number[2];
assign weights[1] = ~random_number[9] & ~random_number[8] & ~random_number[7] & ~random_number[6] & 
				~random_number[5] & ~random_number[4] & ~random_number[3] & 
				~random_number[2] & random_number[1];
assign weights[0] = ~random_number[9] & ~random_number[8] & ~random_number[7] & ~random_number[6] & 
				~random_number[5] & ~random_number[4] & ~random_number[3] & 
				~random_number[2] & ~random_number[1] & random_number[0];

// Calculate intermediate values
for (i = 0; i < 10; i = i + 1) assign intermediates[i] = weights[i] & binary_number[i];

// Use intermediate values to determine the next value in the bitstream
assign stochastic_number = |intermediates;

endmodule
